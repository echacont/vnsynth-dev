// ELeonora Chacón Taylor 2024
// wavetable.vh wavetable hardware description header file

`define WAVE_BRAM_DATA_WIDTH    16
`define WAVE_BRAM_DATA_SIZE     2048
`define WAVE_BRAM_ADDR_WIDTH    11

