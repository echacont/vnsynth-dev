// ELeonora Chacón Taylor 2024
// wavetable_top.v wavetable hardware description top file

`include "wavetable.vh"

module wavetable_top ( 
        input  i_clk, 
        input  i_reset,
		// Wishbone interface
		input  i_wb_cyc, 
        input  i_wb_stb, 
        input         i_wb_we, 
        input  [5:0]  i_wb_addr, 
        input  [31:0] i_wb_data,
		output reg o_wb_ack = 0, 
        output o_wb_stall, 
        output reg [31:0] o_wb_data = 0,
        // Pulse density modulation audio output
		output o_pdm); 

    // Wishbone register write enable
    wire reg_we = i_wb_cyc & i_wb_stb & i_wb_we & !o_wb_ack;
    
    always @(posedge i_clk) begin

        o_wb_ack <= i_wb_cyc & !o_wb_ack; // Always acknowledge
        // these signals need to be only a pulse
        wram_we <= 0;
        wram_en <= 0;
        stop_synth <= 0;
        start_synth <= 0;

        // Wishbone write address decoder
        // FIXME: there is potential bug:
        // it should not be possible to write the RAM while synthesis is on.
        if (reg_we)
            case (i_wb_addr[5:2])
                // wavetable ram control
                0: begin
                    wram_we   <= i_wb_data[0];
                    wram_en   <= 1;
                end
                // wavetable ram address
                // logic was moved below
                //1: wram_addr <= i_wb_data[`WAVE_BRAM_DATA_WIDTH-1:0];
                // wavetable ram data in
                2: wram_di   <= i_wb_data[`WAVE_BRAM_DATA_WIDTH-1:0];
                // synthesis control
                3: begin
                    stop_synth  <= i_wb_data[1];
                    start_synth  <= i_wb_data[0];
                end
                // synthesis wave sample lenght
                4: wram_length <= i_wb_data[11:0];
                // synthesis: pdmaudio reload timer
                5: begin
                   pdm_timer <= i_wb_data[15:0]; 
                end

            endcase

        // Wishbone read address decoder
        if (~reg_we)
            case (i_wb_addr[5:2])
                // status register 
                0: o_wb_data <= 0;
                // wavetable ram address
                1: o_wb_data[`WAVE_BRAM_DATA_WIDTH-1:0] <= wram_addr;
                // wavetable ram data out
                2: o_wb_data[`WAVE_BRAM_DATA_WIDTH-1:0] <= wram_dout;
            endcase
    end

    // Wavetable RAM signals
    wire [`WAVE_BRAM_DATA_WIDTH-1:0]  wram_dout;
    wire [`WAVE_BRAM_ADDR_WIDTH-1:0]  next_wram_addr;
    
    // registers
    reg   wram_we = 0;
    reg   wram_en = 0;
    reg   wram_en_read;
    wire  wram_en_or;
    reg  [`WAVE_BRAM_DATA_WIDTH-1:0]  wram_di = 0;
    reg  [`WAVE_BRAM_ADDR_WIDTH-1:0]  wram_addr = 0;
    reg  [11:0] wram_length = `WAVE_CYCLE_LENGTH;
    reg  inc_wram_addr = 0;
    reg  reset_wram_addr = 0;

    assign next_wram_addr = wram_addr + 1;
    assign wram_en_or = wram_en | wram_en_read;

    // wram address logic
    always @(posedge i_clk) begin
        // wishbone write addressing wram_addr register
        if (reg_we & (i_wb_addr[5:2] == 1)) 
            wram_addr <= i_wb_data[`WAVE_BRAM_DATA_WIDTH-1:0];
        // pdmaudio operation requires the next sample
        else if (inc_wram_addr) begin
            if (next_wram_addr < wram_length) wram_addr <= next_wram_addr;
            else wram_addr <= 0;
        end
        else if (reset_wram_addr) wram_addr <= 0;
        else wram_addr <= wram_addr;
    end

    // BRAM instance
    rams_sp_nc wave_bram0 (
        .clk    (i_clk),
        .we     (wram_we),
        .en     (wram_en_or),
        .addr   (wram_addr),
        .di     (wram_di),
        .dout   (wram_dout));

    // synthesizer state
    reg start_synth = 0;    // signal generated by wishbone write
    reg stop_synth = 1;     // signal generated by wishbone write
    reg audio_en = 0;       // enables the PDM engine
    reg [1:0] synth_state = `SYNTH_FSM_IDLE;
    reg [1:0] next_synth_state = `SYNTH_FSM_IDLE;
    // PDM audio
    reg pdm_reset = 0;
    reg [1:0] pdm_state = `PDM_FSM_IDLE;
    reg [1:0] next_pdm_state = `PDM_FSM_IDLE;
    reg pdm_cyc  = 0;
    reg pdm_we   = 0;
    reg pdm_addr = 0;
    reg [`WAVE_PDM_DATA_WIDTH-1:0] pdm_data = 0;
    reg [15:0] pdm_timer = 16'd1133;
    reg pdm_timer_update = 0;
    wire pdm_reset_w;
    assign pdm_reset_w = i_reset | pdm_reset;

    // main synthesis FSM
    // Enables PDM engine and controls wavetable RAM pointers
    always @(posedge i_clk) begin
        pdm_reset <= 0;
        audio_en <= 0;
        reset_wram_addr <= 0;
        case (synth_state)
            // Idle (no synthesis, silence, off)
            `SYNTH_FSM_IDLE: begin
                if (stop_synth) next_synth_state <= `SYNTH_FSM_IDLE;
                else if (start_synth) next_synth_state <= `SYNTH_FSM_RESET; 
                else next_synth_state <= `SYNTH_FSM_IDLE;
            end
            // reset pdmaudio
            `SYNTH_FSM_RESET: begin
                pdm_reset <= 1;
                next_synth_state <= `SYNTH_FSM_SETUP;
            end
            // setup (reset wram address pointer)
            `SYNTH_FSM_SETUP: begin
                reset_wram_addr <= 1;
                // wait until PDM audio is ready
                if (next_pdm_state == `PDM_FSM_IDLE) 
                    next_synth_state <= `SYNTH_FSM_AUDIO;
                else next_synth_state <= `SYNTH_FSM_SETUP;
            end
            // synthesis/audio on
            `SYNTH_FSM_AUDIO: begin
                audio_en <= 1;
                if (stop_synth) begin
                    next_synth_state <= `SYNTH_FSM_IDLE;
                end
                else next_synth_state <= `SYNTH_FSM_AUDIO;
            end
        endcase
    end

    // PDM audio FSM.
    // Controls operation of PDM audio engine
    always @(posedge i_clk) begin
        wram_en_read <= 0;
        inc_wram_addr <= 0;
        case (pdm_state)
            // Idle
            `PDM_FSM_IDLE: begin
                pdm_cyc  <= 0;
                pdm_we   <= 0;
                pdm_addr <= 0;
                // synth is initializing
                // or pdm engine needs a new sample
                // prepare inputs to reload pwmaudio registers
                // signal read to wave ram using current wram address
                if ((next_synth_state == `SYNTH_FSM_SETUP) | (pdm_int & audio_en)) begin
                    wram_en_read <= 1;
                    next_pdm_state <= `PDM_FSM_READ_SAMPLE;
                end
                // nothing to do
                else next_pdm_state <= `PDM_FSM_IDLE;
            end
            // Read sample from wavetable RAM
            // prepare inputs to pwm audio
            `PDM_FSM_READ_SAMPLE: begin
                // wait until cycle is complete, 
                // move wram read data out to pdm_data bus
                // and prepare inputs to pdmaudio
                if (~wram_en_read) begin
                    pdm_data  <= wram_dout;
                    pdm_cyc   <= 1;
                    pdm_we    <= 1;
                    pdm_addr  <= 0;
                    next_pdm_state <= `PDM_FSM_WRITE_SAMPLE;
                end
            end
            // Write sample
            `PDM_FSM_WRITE_SAMPLE: begin
                // wait until pwmaudio acks 
                // set next wram address
                // if setup, we also need to write reload timer
                if (pdm_ack) begin
                    if ((next_synth_state == `SYNTH_FSM_SETUP) | pdm_timer_update)  begin
                        pdm_cyc  <= 1;
                        pdm_we   <= 1;
                        pdm_addr <= 1;
                        pdm_data <= pdm_timer;
                        next_pdm_state <= `PDM_FSM_WRITE_RELOAD;
                    end
                    // else (only ack) pdmaudio is on
                    // we are done, return PDM FSM to idle
                    else begin
                        pdm_cyc   <= 0;
                        pdm_we    <= 0;
                        next_pdm_state <= `PDM_FSM_IDLE;
                    end
                    inc_wram_addr <= 1;
                end
                else  next_pdm_state <= `PDM_FSM_WRITE_SAMPLE;
            end
            // Write reload value
            `PDM_FSM_WRITE_RELOAD: begin
                // wait until pwmaudio acks to bring down lines
                if (pdm_ack) begin
                    pdm_cyc  <= 0;
                    pdm_we   <= 0;
                    pdm_addr <= 0;
                    wram_en_read  <= 1;
                    next_pdm_state <= `PDM_FSM_IDLE;
                end
                else next_pdm_state <= `PDM_FSM_WRITE_RELOAD;
            end
        endcase     
    end

    always @(negedge i_clk) begin
        synth_state <= next_synth_state; 
        pdm_state <= next_pdm_state; 
    end

    wire [31:0] pdm_data_out;
    wire pdm_ack;

    wire pdm_int;
    wire pdm_clk;

    // gate PDM clock if synth state idle
    assign pdm_clk = i_clk & (synth_state != `SYNTH_FSM_IDLE);

    wbpdmaudio_mod pdmaudio0 (
        .i_clk      (pdm_clk),
        .i_reset    (pdm_reset_w),
        .i_wb_cyc   (pdm_cyc),
        .i_wb_stb   (pdm_cyc),
        .i_wb_we    (pdm_we),
        .i_wb_addr  (pdm_addr),
        .i_wb_data  (pdm_data),
        .o_wb_ack   (pdm_ack),
        .o_wb_data  (pdm_data_out),
        .o_pdm      (o_pdm),
        .o_int      (pdm_int));

endmodule

// elecha: using example code from Xilinx:
// Single-Port Block RAM No-Change Mode
// File: rams_sp_nc.v

module rams_sp_nc (clk, we, en, addr, di, dout);

input clk; 
input we; 
input en;
input [`WAVE_BRAM_ADDR_WIDTH-1:0] addr; 
input [`WAVE_BRAM_DATA_WIDTH-1:0] di; 
output [`WAVE_BRAM_DATA_WIDTH-1:0] dout;

reg [`WAVE_BRAM_DATA_WIDTH-1:0] RAM [`WAVE_BRAM_DATA_SIZE-1:0];
reg [`WAVE_BRAM_DATA_WIDTH-1:0] dout;

always @(posedge clk)
begin
  if (en)
  begin
    if (we)
      RAM[addr] <= di;
    else
      dout <= RAM[addr];
  end
end
endmodule

// reusing code from Dan Gisselquist's wbpwmaudio controller
// with some fixes due to bug related to i_wb_cyc and how data is passed to
// the pulse density modulator, which was itself replaced with 
// other design.
// wishbone interface is emulated by the wavetable logic
module	wbpdmaudio_mod (i_clk, i_reset,
		// Wishbone interface
		i_wb_cyc, i_wb_stb, i_wb_we, i_wb_addr, i_wb_data,
			o_wb_ack, o_wb_stall, o_wb_data,
		o_pdm, o_aux, o_int);
	parameter DEFAULT_RELOAD = 16'd1133,  // about 44.1 kHz @ 50 MHz
            //DEFAULT_RELOAD = 16'd1814, // about 44.1 kHz @  80MHz
			//DEFAULT_RELOAD = 16'd2268,//about 44.1 kHz @ 100MHz
			NAUX=2, // Dev control values
			VARIABLE_RATE=1,
			TIMING_BITS=16;
	input	wire		i_clk, i_reset;
	input	wire		i_wb_cyc, i_wb_stb, i_wb_we;
	input	wire		i_wb_addr;
	input	wire	[31:0]	i_wb_data;
	output	reg		o_wb_ack;
	output	wire		o_wb_stall;
	output	wire	[31:0]	o_wb_data;
	output	wire		o_pdm;
	output	reg	[(NAUX-1):0]	o_aux;
	output	wire		o_int;


	// How often shall we create an interrupt?  Every reload_value clocks!
	// If VARIABLE_RATE==0, this value will never change and will be kept
	// at the default reload rate (defined up top)
	wire	[(TIMING_BITS-1):0]	w_reload_value;
	generate
	if (VARIABLE_RATE != 0)
	begin
		reg	[(TIMING_BITS-1):0]	r_reload_value;
		initial	r_reload_value = DEFAULT_RELOAD;
		always @(posedge i_clk) // Data write
            // Eleonora Chacon: adding i_wb_cyc to this condition
			if ((i_wb_cyc)&&(i_wb_stb)&&(i_wb_addr)&&(i_wb_we))
				r_reload_value <= i_wb_data[(TIMING_BITS-1):0] - 1'b1;
		assign	w_reload_value = r_reload_value;
	end else begin
		assign	w_reload_value = DEFAULT_RELOAD;
	end endgenerate

	//
	// The next value timer
	//
	// We'll want a new sample every w_reload_value clocks.  When the
	// timer hits zero, the signal ztimer (zero timer) will also be
	// set--allowing following logic to depend upon it.
	//
	reg				ztimer;
	reg	[(TIMING_BITS-1):0]	timer;
	initial	timer = DEFAULT_RELOAD;
	initial	ztimer= 1'b0;
	always @(posedge i_clk)
		if (i_reset)
			ztimer <= 1'b0;
		else
			ztimer <= (timer == { {(TIMING_BITS-1){1'b0}}, 1'b1 });

	always @(posedge i_clk)
		if ((ztimer)||(i_reset))
			timer <= w_reload_value;
		else
			timer <= timer - {{(TIMING_BITS-1){1'b0}},1'b1};

	//
	// Whenever the timer runs out, accept the next value from the single
	// sample buffer.
	//
	reg	[15:0]	sample_out;
	always @(posedge i_clk)
		if (ztimer)
			sample_out <= next_sample;

	//
	// Control what's in the single sample buffer, next_sample, as well as
	// whether or not it's a valid sample.  Specifically, if next_valid is
	// false, then the sample buffer needs a new value.  Once the buffer
	// has a value within it, further writes will just quietly overwrite
	// this value.
	reg	[15:0]	next_sample;
	reg		next_valid;
	initial	next_valid = 1'b1;
	initial	next_sample = 16'h8000;
	always @(posedge i_clk) // Data write
        // Eleonora Chacon: adding i_wb_cyc to this condition
		if ((i_wb_stb)&&(i_wb_we)&&(i_wb_cyc)
				&&((!i_wb_addr)||(VARIABLE_RATE==0)))
		begin
			// Write with two's complement data, convert it
			// internally to an unsigned binary offset
			// representation
            next_sample <= { !i_wb_data[15], i_wb_data[14:0] };
			next_valid <= 1'b1;
		end else if (ztimer)
			next_valid <= 1'b0;

	// If the value in our sample buffer isn't valid, create an interrupt
	// that can be sent to a processor to know when to send a new sample.
	// This output can also be used to control a read from a FIFO as well,
	// depending on how you wish to use the core.
	assign	o_int = (!next_valid);

    // Eleonora Chacon
    // To generate our waveform, I will use a different PDM method

    wire pdm_out;

    pdm pdm0(
        .clk    (i_clk),
        .rst    (i_reset),
        .din    (sample_out),
        .dout   (pdm_out),
        .error  ());

    //assign o_pdm = ~pdm_out ? 1'b0 : 1'bz;
    assign o_pdm = pdm_out;

	// Handle the bus return traffic.
	generate
	if (VARIABLE_RATE == 0)
	begin
		// If we are running off of a fixed rate, then just return
		// the current setting of the aux registers, the current
		// interrupt value, and the current sample we are outputting.
		assign o_wb_data = { {(12-NAUX){1'b0}}, o_aux,
					3'h0, o_int, sample_out };
	end else begin
		// On the other hand, if we have been built to support a
		// variable sample rate, then return the reload value for
		// address one but otherwise the data value (above) for address
		// zero.
		reg	[31:0]	r_wb_data;
		always @(posedge i_clk)
			if (i_wb_addr)
				r_wb_data <= { (32-TIMING_BITS),w_reload_value};
			else
				r_wb_data <= { {(12-NAUX){1'b0}}, o_aux,
						3'h0, o_int, sample_out };
		assign	o_wb_data = r_wb_data;
	end endgenerate

	// Always ack on the clock following any request
	initial	o_wb_ack = 1'b0;
	always @(posedge i_clk)
		o_wb_ack <= (i_wb_stb);

	// Never stall
	assign	o_wb_stall = 1'b0;

	// Make Verilator happy.  Since we aren't using all of the bits from
	// the bus, Verilator -Wall will complain.  This just informs
	// V*rilator that we already know these bits aren't being used.
	//
	// verilator lint_off UNUSED
	wire	[14:0] unused;
	assign	unused = {i_wb_data[31:21], i_wb_data[19:17] };
	// verilator lint_on  UNUSED

endmodule

// Pulse Density Modulation code taken from
// https://www.koheron.com/blog/2016/09/27/pulse-density-modulation
module pdm #(parameter NBITS = 16)
(
  input wire                      clk,
  input wire [NBITS-1:0]          din,
  input wire                      rst,
  output reg                      dout,
  output reg [NBITS-1:0]          error
);

  localparam integer MAX = 2**NBITS - 1;
  reg [NBITS-1:0] din_reg;
  reg [NBITS-1:0] error_0;
  reg [NBITS-1:0] error_1;

  always @(posedge clk) begin
    din_reg <= din;
    error_1 <= error + MAX - din_reg;
    error_0 <= error - din_reg;
  end

  always @(posedge clk) begin
    if (rst == 1'b1) begin
      dout <= 0;
      error <= 0;
    end
    else if (din_reg >= error) begin
      dout <= 1;
      error <= error_1;
    end else begin
      dout <= 0;
      error <= error_0;
    end
  end

endmodule
